/*
   Copyright 2024 jackkyyang

   Licensed under the Apache License, Version 2.0 (the "License");
   you may not use this file except in compliance with the License.
   You may obtain a copy of the License at

       http://www.apache.org/licenses/LICENSE-2.0

   Unless required by applicable law or agreed to in writing, software
   distributed under the License is distributed on an "AS IS" BASIS,
   WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
   See the License for the specific language governing permissions and
   limitations under the License.

 ***************************************************************************
 * File Name: cmprs_4to2.sv
 * Creation Date: 2024/10/20
 * Author: jackkyyang
 * Description:
 *  a fast 4-to-2 compressor.
 *  the weight of each output is the weight of input + 1
 ***************************************************************************
*/

module cmprs_4to2
#(
    parameter integer WIDTH = 1
)
(
    input  logic [WIDTH-1:0] cin,     // carry in
    input  logic [WIDTH-1:0] a,       // input a
    input  logic [WIDTH-1:0] b,       // input b
    input  logic [WIDTH-1:0] c,       // input c
    input  logic [WIDTH-1:0] d,       // input d
    output logic [WIDTH-1:0] cout_a,  // carry out
    output logic [WIDTH-1:0] cout_b,  // carry out
    output logic [WIDTH-1:0] sum      // sum
);

  wire[WIDTH-1:0] xor_ab = a ^ b;
  wire[WIDTH-1:0] xor_cd = c ^ d;

  wire[WIDTH-1:0] xor_abcd = (xor_ab ^ xor_cd);

  assign sum = xor_abcd ^ cin;
  assign cout_a = (xor_abcd & cin) | ((~xor_abcd) & d);
  assign cout_b = (a & b) | (b & c) | (a & c);


endmodule
